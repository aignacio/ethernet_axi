`ifndef _UTILS_PKG_
`define _UTILS_PKG_
  package utils_pkg;
    `include "axi_pkg.svh"
    `include "eth_pkg.svh"
  endpackage
`endif
