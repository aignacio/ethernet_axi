/**
 * File              : axi_bridge.sv
 * License           : MIT license <Check LICENSE>
 * Author            : Anderson Ignacio da Silva (aignacio) <anderson@aignacio.com>
 * Date              : 19.07.2022
 * Last Modified Date: 19.07.2022
 */

